module top(

);

endmodule
